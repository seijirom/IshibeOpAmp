* Created by KLayout

* cell 1umiv
.SUBCKT 1umiv
* net 1 Vdd
* net 2 Vout
* net 4 VINM
* net 5 VINP
* net 6 SUBSTRATE
* device instance $1 r0 *1 102.5,72 CAP
C$1 2 3 2.9952e-12
* device instance $2 r0 *1 5.5,141 HRES
R$2 7 1 40250
* device instance $3 m90 *1 72,63 NMOS
M$3 6 8 2 6 NMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $4 m90 *1 72,99 NMOS
M$4 6 8 2 6 NMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $5 r0 *1 65.5,63 NMOS
M$5 6 8 2 6 NMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $6 r0 *1 65.5,99 NMOS
M$6 6 8 2 6 NMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $7 r0 *1 24,24.5 NMOS
M$7 6 7 12 6 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $8 r0 *1 12.5,24.5 NMOS
M$8 6 7 7 6 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $9 m90 *1 66.5,31.5 NMOS
M$9 8 3 1 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $10 r0 *1 52.5,15.5 NMOS
M$10 6 14 8 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $11 r0 *1 46,42 NMOS
M$11 17 9 3 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $12 m90 *1 39.5,42 NMOS
M$12 14 9 9 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $13 m45 *1 16,53.5 NMOS
M$13 6 7 15 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $14 r0 *1 39.5,15.5 NMOS
M$14 6 14 14 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $15 m90 *1 46,15.5 NMOS
M$15 6 14 17 6 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $16 m90 *1 50.5,69 PMOS
M$16 10 15 3 10 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $17 r0 *1 36,69 PMOS
M$17 11 15 9 11 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $18 r0 *1 12.5,104.5 PMOS
M$18 16 13 13 16 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $19 m90 *1 21.5,104.5 PMOS
M$19 16 13 13 16 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $20 m90 *1 21.5,73.5 PMOS
M$20 13 15 15 13 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $21 r0 *1 12.5,73.5 PMOS
M$21 13 15 15 13 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $22 m90 *1 48.5,101.5 PMOS
M$22 16 4 10 16 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $23 r0 *1 39.5,101.5 PMOS
M$23 16 5 11 16 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $24 m90 *1 23.5,139 PMOS
M$24 1 12 12 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $25 r0 *1 14.5,139 PMOS
M$25 1 12 12 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $26 m90 *1 73,139 PMOS
M$26 1 12 2 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $27 m90 *1 48.5,139 PMOS
M$27 1 12 16 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $28 r0 *1 39.5,139 PMOS
M$28 1 12 16 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $29 r0 *1 64,139 PMOS
M$29 1 12 2 1 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
.ENDS 1umiv
