* Created by KLayout

* cell 1umiv
.SUBCKT 1umiv
* net 2 Vdd
* net 5 Vbias
* net 9 VINM
* net 11 Vout
* net 12 VINP
* net 17 Gnd
* device instance $1 r0 *1 23,139 PMOS
M$1 2 10 10 2 PMOS L=1U W=50U AS=100P AD=100P PS=83U PD=83U
* device instance $3 r0 *1 48.5,101.5 PMOS
M$3 7 9 15 15 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $4 r0 *1 48.5,139 PMOS
M$4 15 10 2 2 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $5 r0 *1 73,139 PMOS
M$5 11 10 2 2 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $8 r0 *1 39.5,101.5 PMOS
M$8 15 12 6 15 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $9 r180 *1 11.5,141.5 HRES
R$9 2 5 40250 HRES
* device instance $10 m90 *1 72.5,68.5 NMOS
M$10 17 3 11 17 NMOS L=1U W=100U AS=200P AD=200P PS=216U PD=216U
* device instance $14 r0 *1 12.5,23 NMOS
M$14 17 5 5 17 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $15 r0 *1 24,23 NMOS
M$15 17 5 10 17 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $16 m90 *1 59,37.5 NMOS
M$16 3 4 2 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $17 r0 *1 53,14 NMOS
M$17 17 13 3 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $18 r0 *1 46,40.5 NMOS
M$18 16 8 4 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $19 m45 *1 16,52 NMOS
M$19 17 5 14 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $20 m90 *1 39,40.5 NMOS
M$20 13 8 8 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $21 m90 *1 46,14 NMOS
M$21 17 13 16 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $22 r0 *1 39,14 NMOS
M$22 17 13 13 17 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $23 r0 *1 12.5,104.5 PMOS
M$23 15 1 1 15 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $24 r0 *1 12.5,73.5 PMOS
M$24 1 14 14 1 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $27 m90 *1 50.5,67.5 PMOS
M$27 7 14 4 7 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $28 r0 *1 36,67.5 PMOS
M$28 6 14 8 6 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $29 m90 *1 82,22.5 CAP
C$29 11 4 3.0186e-12 CAP
.ENDS 1umiv
