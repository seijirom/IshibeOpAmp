* Created by KLayout

* cell 1umiv
.SUBCKT 1umiv
* net 1 Vbias
* net 2 Vdd
* net 4 Vout
* net 5 VINM
* net 6 VINP
* net 7 Gnd
* device instance $1 r0 *1 102.5,72 CAP
C$1 4 3 2.9952e-12
* device instance $2 r0 *1 2,141 HRES
R$2 1 2 40250
* device instance $3 m90 *1 72.5,61.5 NMOS
M$3 7 8 4 7 NMOS L=1U W=100U AS=200P AD=200P PS=216U PD=216U
* device instance $7 r0 *1 12.5,23 NMOS
M$7 7 1 1 7 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $8 r0 *1 24,23 NMOS
M$8 7 1 13 7 NMOS L=1U W=34U AS=68P AD=68P PS=72U PD=72U
* device instance $9 m90 *1 66.5,30 NMOS
M$9 8 3 2 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $10 r0 *1 53,14 NMOS
M$10 7 14 8 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $11 r0 *1 46,40.5 NMOS
M$11 17 9 3 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $12 m90 *1 39,40.5 NMOS
M$12 14 9 9 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $13 m45 *1 16,52 NMOS
M$13 7 1 15 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $14 r0 *1 39,14 NMOS
M$14 7 14 14 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $15 m90 *1 46,14 NMOS
M$15 7 14 17 7 NMOS L=1U W=16U AS=32P AD=32P PS=36U PD=36U
* device instance $16 m90 *1 50.5,67.5 PMOS
M$16 10 15 3 10 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $17 r0 *1 36,67.5 PMOS
M$17 11 15 9 11 PMOS L=1U W=19U AS=38P AD=38P PS=42U PD=42U
* device instance $18 r0 *1 12.5,104.5 PMOS
M$18 16 12 12 16 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $20 m90 *1 21.5,73.5 PMOS
M$20 12 15 15 12 PMOS L=1U W=38U AS=76P AD=76P PS=84U PD=84U
* device instance $22 m90 *1 48.5,101.5 PMOS
M$22 16 5 10 16 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $23 r0 *1 39.5,101.5 PMOS
M$23 16 6 11 16 PMOS L=1U W=25U AS=50P AD=50P PS=54U PD=54U
* device instance $24 m90 *1 23.5,139 PMOS
M$24 2 13 13 2 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $25 m90 *1 48.5,139 PMOS
M$25 2 13 16 2 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
* device instance $26 m90 *1 73,139 PMOS
M$26 2 13 4 2 PMOS L=1U W=50U AS=100P AD=100P PS=108U PD=108U
.ENDS 1umiv
