* Z:\HOME\SEIJIROM\WORK\2021_9\ISHIBEOPAMP\ISHIBE_TB.ASC
*XX1 N004 N001 OUT N002 NC_01 OPAMP3UREIAUTO
*R1 N004 N003 10K
*R2 OUT N004 100K
*V1 N003 N001 SINE(0 0.1 1K) AC 1
*V2 N002 N001 3
*V3 N001 0 3
*
* BLOCK SYMBOL DEFINITIONS
.SUBCKT OPAMP3UREIAUTO VINM VINP VOUT VDD VBIAS
M1 N010 N010 0 0 NMOS L=1U W=16U
M2 N008 N008 N010 0 NMOS L=1U W=16U
M3 N011 N010 0 0 NMOS L=1U W=16U
M4 N007 N008 N011 0 NMOS L=1U W=16U
M5 N001 VBIAS 0 0 NMOS L=1U W=34U
M6 N006 VBIAS 0 0 NMOS L=1U W=16U
M10 VOUT N009 0 0 NMOS L=1U W=100U
M11 N009 N010 0 0 NMOS L=1U W=16U
M12 VDD N007 N009 0 NMOS L=1U W=16U
M13 N002 N001 VDD VDD PMOS L=1U W=50U
M14 N003 N003 N002 N002 PMOS L=1U W=38U
M15 N006 N006 N003 N003 PMOS L=1U W=38U
M16 N007 N006 N005 N005 PMOS L=1U W=19U
M17 N008 N006 N004 N004 PMOS L=1U W=19U
M18 N004 VINM N002 N002 PMOS L=1U W=25U
M20 VOUT N001 VDD VDD PMOS L=1U W=50U
M21 N005 VINP N002 N002 PMOS L=1U W=25U
M24 N001 N001 VDD VDD PMOS L=1U W=50U
M7 VBIAS VBIAS 0 0 NMOS L=1U W=34U
R1 VDD VBIAS 40K
C1 VOUT N007 3P
*.INC ./MODELS/OR1_MOS
*.INCLUDE "./BSIM3V3N.MOD"
*.INCLUDE "./BSIM3V3P.MOD"
.ENDS OPAMP3UREIAUTO

.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\SEIJIROM\DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
*.INCLUDE MODELS/OR1_MOS
*.INCLUDE "./BSIM3V3N.MOD"
*.INCLUDE "./BSIM3V3P.MOD"
.AC DEC 10 1 1G
.BACKANNO
.GLOBAL 0
.END
