* Z:\HOME\ANAGIX\ALBDATA\4802\1UMTESTBE.ASC
*XX1 NC_01 NC_02 N001 N005 N002 N002 1UMCONTROL
*XX2 NC_03 N001 N004 N002 N003 N003 1UMIV_CONV
*V1 N005 0 2.5
*V2 N001 0 5
*V3 N004 0 2.5
*
* BLOCK SYMBOL DEFINITIONS
*.SUBCKT 1UMCONTROL VBIAS_CE VBIAS_RE VDD VIN CE RE
*XX1 N001 RE N001 VDD VBIAS_RE OPAMP3UREIAUTO
*XX2 N001 VIN CE VDD VBIAS_CE OPAMP3UREIAUTO
*.ENDS 1UMCONTROL
*
*.SUBCKT 1UMIV_CONV VBIAS_WE VDD VDD_HALF WE R1K VOUT
*XX1 WE VDD_HALF VOUT VDD VBIAS_WE OPAMP3UREIAUTO
*R1 R1K WE 1K
*.ENDS 1UMIV_CONV
*
.SUBCKT OPAMP3UREIAUTO VINM VINP VOUT VDD VBIAS
M1 N010 N010 0 0 NMOS L=1U W=16U
M2 N008 N008 N010 0 NMOS L=1U W=16U
M3 N011 N010 0 0 NMOS L=1U W=16U
M4 N007 N008 N011 0 NMOS L=1U W=16U
M5 N001 VBIAS 0 0 NMOS L=1U W=34U
M6 N006 VBIAS 0 0 NMOS L=1U W=16U
M10 VOUT N009 0 0 NMOS L=1U W=100U
M11 N009 N010 0 0 NMOS L=1U W=16U
M12 VDD N007 N009 0 NMOS L=1U W=16U
M13 N002 N001 VDD VDD PMOS L=1U W=50U
M14 N003 N003 N002 N002 PMOS L=1U W=38U
M15 N006 N006 N003 N003 PMOS L=1U W=38U
M16 N007 N006 N005 N005 PMOS L=1U W=19U
M17 N008 N006 N004 N004 PMOS L=1U W=19U
M18 N004 VINM N002 N002 PMOS L=1U W=25U
M20 VOUT N001 VDD VDD PMOS L=1U W=50U
M21 N005 VINP N002 N002 PMOS L=1U W=25U
M24 N001 N001 VDD VDD PMOS L=1U W=50U
M7 VBIAS VBIAS 0 0 NMOS L=1U W=34U
R1 VDD VBIAS 40K
C1 VOUT N007 3P
*.INC ./MODELS/OR1_MOS
*.INCLUDE "./BSIM3V3N.MOD"
*.INCLUDE "./BSIM3V3P.MOD"
.ENDS OPAMP3UREIAUTO

.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\ANAGIX\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
.MODEL NMOS NMOS
.MODEL PMOS PMOS
*.INCLUDE "./MODELS/OR1_MOS"
.OP
.BACKANNO
.BACKANNO
.END
