.TITLE KICAD SCHEMATIC
M11 NET__M10_PAD3_ NET__M10_PAD3_ "/GND" "/GND" NMOS L=1U W=16U
M10 NET__M10_PAD1_ NET__M10_PAD1_ NET__M10_PAD3_ "/GND" NMOS L=1U W=16U
M14 NET__M13_PAD3_ NET__M10_PAD3_ "/GND" "/GND" NMOS L=1U W=16U
M13 NET__C1_PAD2_ NET__M10_PAD1_ NET__M13_PAD3_ "/GND" NMOS L=1U W=16U
M2 NET__M18_PAD2_ NET__M1_PAD1_ "/GND" "/GND" NMOS L=1U W=34U
M4 NET__M12_PAD2_ NET__M1_PAD1_ "/GND" "/GND" NMOS L=1U W=16U
M19 "/VOUT" NET__M16_PAD3_ "/GND" "/GND" NMOS L=1U W=100U
M17 NET__M16_PAD3_ NET__M10_PAD3_ "/GND" "/GND" NMOS L=1U W=16U
M16 "/VDD" NET__C1_PAD2_ NET__M16_PAD3_ "/GND" NMOS L=1U W=16U
M8 NET__M15_PAD3_ NET__M18_PAD2_ "/VDD" "/VDD" PMOS L=1U W=50U
M5 NET__M5_PAD1_ NET__M5_PAD1_ NET__M15_PAD3_ NET__M15_PAD3_ PMOS L=1U W=38U
M6 NET__M12_PAD2_ NET__M12_PAD2_ NET__M5_PAD1_ NET__M5_PAD1_ PMOS L=1U W=38U
M12 NET__C1_PAD2_ NET__M12_PAD2_ NET__M12_PAD3_ NET__M12_PAD3_ PMOS L=1U W=19U
M9 NET__M10_PAD1_ NET__M12_PAD2_ NET__M7_PAD1_ NET__M7_PAD1_ PMOS L=1U W=19U
M7 NET__M7_PAD1_ NC_01 NET__M15_PAD3_ NET__M15_PAD3_ PMOS L=1U W=25U
M18 "/VOUT" NET__M18_PAD2_ "/VDD" "/VDD" PMOS L=1U W=50U
M3 NET__M18_PAD2_ NET__M18_PAD2_ "/VDD" "/VDD" PMOS L=1U W=50U
M1 NET__M1_PAD1_ NET__M1_PAD1_ "/GND" "/GND" NMOS L=1U W=34U
R3 "/VDD" NET__M1_PAD1_ 40K
C1 "/VOUT" NET__C1_PAD2_ 3P
M15 NET__M12_PAD3_ NC_02 NET__M15_PAD3_ NET__M15_PAD3_ PMOS L=1U W=25U
.END
